`include "fifo_pkg.sv"
`include "fifo_trans.sv"
`include "fifo_if.sv"
`include "fifo_sequencer.sv"
`include "fifo_monitor.sv"
`include "fifo_fcov.sv"
`include "fifo_scoreboard.sv"
`include "fifo_dri.sv"
`include "fifo_agent.sv"
`include "fifo_env.sv"
`include "fifo_sequence.sv"
`include "fifo_base_test.sv"
`include "fifo_rand_test.sv"
